module decoder_tb();

  logic        clk;
  logic        reset_n;
  logic        ID;
  logic [31:0] i_data_read;

  logic d_write_enable;
  logic d_load_enable;
  logic Iv_alu;
  logic Pc_alu;
  logic [1:0] Pc_cmd;
  logic [1:0] Pc_val;
  logic [3:0] I;
  logic [4:0] Rs1;
  logic [4:0] Rs2;
  logic [4:0] Rd;
  logic [31:0] Iv;

  always
    begin
      #5ns
      clk <= !clk;
    end

  initial
    begin
      #1ns
      clk <= 0;
      reset_n <= 0;
      ID      <= 1;
      #12ns
      reset_n <= 1;

      // On commence par les instructions R
      #10ns
      i_data_read <= 32'b000000,01101,11000,00110,00000,100000;
      #10ns
      i_data_read <= 32'b000000,01101,11000,00110,00000,100100;
      #10ns
      i_data_read <= 32'b000000,01101,11000,00110,00000,100101;
      #10ns
      i_data_read <= 32'b000000,01101,11000,00110,00000,101000;
      #10ns
      i_data_read <= 32'b000000,01101,11000,00110,00000,101100;
      #10ns
      i_data_read <= 32'b000000,01101,11000,00110,00000,000100;
      #10ns
      i_data_read <= 32'b000000,01101,11000,00110,00000,101111;
      #10ns
      i_data_read <= 32'b000000,01101,11000,00110,00000,101001;
      #10ns
      i_data_read <= 32'b000000,01101,11000,00110,00000,000111;
      #10ns
      i_data_read <= 32'b000000,01101,11000,00110,00000,000110;
      #10ns
      i_data_read <= 32'b000000,01101,11000,00110,00000,100010;
      #10ns
      i_data_read <= 32'b000000,01101,11000,00110,00000,100110;

      // Ensuite les deux instructions J
      #10ns
      i_data_read <= 32'b000010,01101110000011000000100110;
      #10ns
      i_data_read <= 32'b000011,01101110000011000000100110;

      // Et enfin les instructions I

      #10ns
      i_data_read <= 32'b001000,01101,11000,0011000000100110;
      #10ns
      i_data_read <= 32'b001100,01101,11000,0011000000100110;
      #10ns
      i_data_read <= 32'b000100,01101,11000,0011000000100110;
      #10ns
      i_data_read <= 32'b000101,01101,11000,0011000000100110;
      #10ns
      i_data_read <= 32'b010011,01101,11000,0011000000100110;
      #10ns
      i_data_read <= 32'b010010,01101,11000,0011000000100110;
      #10ns
      i_data_read <= 32'b001111,01101,11000,0011000000100110;
      #10ns
      i_data_read <= 32'b100011,01101,11000,0011000000100110;
      #10ns
      i_data_read <= 32'b001101,01101,11000,0011000000100110;
      #10ns
      i_data_read <= 32'b011000,01101,11000,0011000000100110;
      #10ns
      i_data_read <= 32'b011100,01101,11000,0011000000100110;
      #10ns
      i_data_read <= 32'b010100,01101,11000,0011000000100110;
      #10ns
      i_data_read <= 32'b011010,01101,11000,0011000000100110;
      #10ns
      i_data_read <= 32'b011001,01101,11000,0011000000100110;
      #10ns
      i_data_read <= 32'b010111,01101,11000,0011000000100110;
      #10ns
      i_data_read <= 32'b010110,01101,11000,0011000000100110;
      #10ns
      i_data_read <= 32'b001010,01101,11000,0011000000100110;
      #10ns
      i_data_read <= 32'b101011,01101,11000,0011000000100110;
      #10ns
      i_data_read <= 32'b001110,01101,11000,0011000000100110;


    end
