module decoder_tb();

  
